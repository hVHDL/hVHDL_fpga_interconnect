library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;

package fpga_interconnect_pkg is

end package fpga_interconnect_pkg;

package body fpga_interconnect_pkg is

end package body fpga_interconnect_pkg;
